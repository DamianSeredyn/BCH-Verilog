module BCH_decoder (

    input  logic        rst,
    input  logic        clk,

   );

    always_ff @(posedge clk or posedge rst)
    begin
	if (rst == 1'b1) 
    begin
        
	end
    else begin
    
    end
end

endmodule