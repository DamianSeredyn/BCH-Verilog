package unit_test_pkg;
    `include "axi4_lite_driver_slave.svh"
endpackage